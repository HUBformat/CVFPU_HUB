// Copyright 2019 ETH Zurich and University of Bologna.
//
// Copyright and related rights are licensed under the Solderpad Hardware
// License, Version 0.51 (the "License"); you may not use this file except in
// compliance with the License. You may obtain a copy of the License at
// http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
// or agreed to in writing, software, hardware and materials distributed under
// this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
// CONDITIONS OF ANY KIND, either express or implied. See the License for the
// specific language governing permissions and limitations under the License.
//
// SPDX-License-Identifier: SHL-0.51

// Author: Stefan Mach <smach@iis.ee.ethz.ch>

module fpnew_opgroup_fmt_slice #(
  parameter fpnew_pkg::opgroup_e     OpGroup       = fpnew_pkg::ADDMUL,
  parameter fpnew_pkg::fp_format_e   FpFormat      = fpnew_pkg::fp_format_e'(0),
  // FPU configuration
  parameter int unsigned             Width         = 32,
  parameter logic                    EnableVectors = 1'b1,
  parameter int unsigned             NumPipeRegs   = 0,
  parameter fpnew_pkg::pipe_config_t PipeConfig    = fpnew_pkg::BEFORE,
  parameter logic                    ExtRegEna     = 1'b0,
  parameter type                     TagType       = logic,
  parameter int unsigned             TrueSIMDClass = 0,
  // Do not change
  localparam int unsigned NUM_OPERANDS = fpnew_pkg::num_operands(OpGroup),
  localparam int unsigned NUM_LANES    = fpnew_pkg::num_lanes(Width, FpFormat, EnableVectors),
  localparam type         MaskType     = logic [NUM_LANES-1:0],
  localparam int unsigned ExtRegEnaWidth = NumPipeRegs == 0 ? 1 : NumPipeRegs
) (
  input logic                               clk_i,
  input logic                               rst_ni,
  // Input signals
  input logic [NUM_OPERANDS-1:0][Width-1:0] operands_i,
  input logic [NUM_OPERANDS-1:0]            is_boxed_i,
  input fpnew_pkg::roundmode_e              rnd_mode_i,
  input fpnew_pkg::operation_e              op_i,
  input logic                               op_mod_i,
  input logic                               vectorial_op_i,
  input TagType                             tag_i,
  input MaskType                            simd_mask_i,
  // Input Handshake
  input  logic                              in_valid_i,
  output logic                              in_ready_o,
  input  logic                              flush_i,
  // Output signals
  output logic [Width-1:0]                  result_o,
  output fpnew_pkg::status_t                status_o,
  output logic                              extension_bit_o,
  output TagType                            tag_o,
  // Output handshake
  output logic                              out_valid_o,
  input  logic                              out_ready_i,
  // Indication of valid data in flight
  output logic                              busy_o,
  // External register enable override
  input  logic [ExtRegEnaWidth-1:0]         reg_ena_i
);

  localparam int unsigned FP_WIDTH  = fpnew_pkg::fp_width(FpFormat);
  localparam int unsigned SIMD_WIDTH = unsigned'(Width/NUM_LANES);


  logic [NUM_LANES-1:0] lane_in_ready, lane_out_valid; // Handshake signals for the lanes
  logic                 vectorial_op;

  logic [NUM_LANES*FP_WIDTH-1:0] slice_result;
  logic [Width-1:0]              slice_regular_result, slice_class_result, slice_vec_class_result;

  fpnew_pkg::status_t    [NUM_LANES-1:0] lane_status;
  logic                  [NUM_LANES-1:0] lane_ext_bit; // only the first one is actually used
  fpnew_pkg::classmask_e [NUM_LANES-1:0] lane_class_mask;
  TagType                [NUM_LANES-1:0] lane_tags; // only the first one is actually used
  logic                  [NUM_LANES-1:0] lane_masks;
  logic                  [NUM_LANES-1:0] lane_vectorial, lane_busy, lane_is_class; // dito

  logic result_is_vector, result_is_class;

  // -----------
  // Input Side
  // -----------
  assign in_ready_o   = lane_in_ready[0]; // Upstream ready is given by first lane
  assign vectorial_op = vectorial_op_i & EnableVectors; // only do vectorial stuff if enabled

  // ---------------
  // Generate Lanes
  // ---------------
  for (genvar lane = 0; lane < int'(NUM_LANES); lane++) begin : gen_num_lanes
    logic [FP_WIDTH-1:0] local_result; // lane-local results
    logic                local_sign;

    // Generate instances only if needed, lane 0 always generated
    if ((lane == 0) || EnableVectors) begin : active_lane
      logic in_valid, out_valid, out_valid_adder, out_valid_mult, out_ready; // lane-local handshake

      logic [NUM_OPERANDS-1:0][FP_WIDTH-1:0] local_operands; // lane-local operands
      logic [FP_WIDTH-1:0]                   op_result;      // lane-local results
      fpnew_pkg::status_t                    op_status;

      assign in_valid = in_valid_i & ((lane == 0) | vectorial_op); // upper lanes only for vectors
      // Slice out the operands for this lane
      always_comb begin : prepare_input
        for (int i = 0; i < int'(NUM_OPERANDS); i++) begin
          local_operands[i] = operands_i[i][(unsigned'(lane)+1)*FP_WIDTH-1:unsigned'(lane)*FP_WIDTH];
        end
      end

      // Instantiate the operation from the selected opgroup
      if (OpGroup == fpnew_pkg::ADDMUL) begin : lane_instance
        
        logic [FP_WIDTH-1:0]  add_result, mult_result;      // lane-local results
        fpnew_pkg::status_t   add_status, mult_status;
        logic                 adder_in_ready, mult_in_ready;
        logic                 adder_out_valid, mult_out_valid;

        fpnew_hub_adder_wrapper #(
          .FpFormat(FpFormat)
        ) i_hub_adder_wrapper (
          .clk_i,
          .rst_ni,
          .operands_i(local_operands),
          .op_i,
          .op_mod_i,
          .in_valid_i(in_valid),
          .in_ready_o(adder_in_ready),
          .flush_i,
          .result_o(add_result),
          .status_o(add_status),
          .out_valid_o(adder_out_valid),
          .out_ready_i(out_ready)
        );
        
        fpnew_hub_multiplier_wrapper #(
          .FpFormat(FpFormat)
        ) i_hub_multiplier_wrapper (
          .clk_i,
          .rst_ni,
          .operands_i(local_operands),
          .op_i,
          .op_mod_i,
          .in_valid_i(in_valid),
          .in_ready_o(mult_in_ready),
          .flush_i,
          .result_o(mult_result),
          .status_o(mult_status),
          .out_valid_o(mult_out_valid),
          .out_ready_i(out_ready)
        );

        // MUX para seleccionar la señal in_ready y las salidas del módulo correcto.
        always_comb begin
          case(op_i)
            fpnew_pkg::ADD: begin
              op_result = add_result;
              op_status = add_status;
              out_valid = adder_out_valid;
              lane_in_ready[lane] = adder_in_ready;
              lane_busy[lane] = 1'b0;
            end
            fpnew_pkg::MUL: begin
              op_result = mult_result;
              op_status = mult_status;
              out_valid = mult_out_valid;
              lane_in_ready[lane] = mult_in_ready;
              lane_busy[lane] = 1'b0;
            end
            default: begin
              op_result = '{default: 1'bx};
              op_status = '{default: 1'bx};
              out_valid = 1'b0;
              lane_in_ready[lane] = 1'b0;
              lane_busy[lane] = 1'b0;
            end
          endcase
        end
        assign lane_is_class[lane]   = 1'b0;
        assign lane_class_mask[lane] = fpnew_pkg::NEGINF;

      end else if (OpGroup == fpnew_pkg::DIVSQRT) begin : lane_instance

        logic [FP_WIDTH-1:0]  div_result, sqrt_result;
        fpnew_pkg::status_t   div_status, sqrt_status;
        logic                 div_in_ready_o, sqrt_in_ready_o;
        logic                 div_start_i, sqrt_start_i;
        logic                 div_out_valid, sqrt_out_valid;
        logic                 div_busy_o, sqrt_busy_o, divsqrt_busy;

        // Instancia del divisor en formato HUB
        fpnew_hub_divider_wrapper #(
          .FpFormat(FpFormat)
        ) i_hub_divider_wrapper (
          .clk_i,
          .rst_ni,
          .operands_i(local_operands), 
          .op_i,
          .op_mod_i,
          .in_valid_i(in_valid),
          .in_ready_o(div_in_ready_o),
          .flush_i,
          .result_o(div_result),
          .status_o(div_status),
          .out_valid_o(div_out_valid),
          .out_ready_i(out_ready),
          .busy_o(div_busy_o)
        );

        fpnew_hub_sqrt_wrapper #(
          .FpFormat(FpFormat)
        ) i_hub_sqrt_wrapper(
          .clk_i(clk_i),
          .rst_ni(rst_ni),
          .operands_i(local_operands),
          .op_i(op_i),
          .op_mod_i(op_mod_i),
          .in_valid_i(in_valid),
          .in_ready_o(sqrt_in_ready_o),
          .flush_i(flush_i),
          .result_o(sqrt_result),
          .status_o(sqrt_status),
          .out_valid_o(sqrt_out_valid),
          .out_ready_i(out_ready),
          .busy_o(sqrt_busy_o)
        );

        // Se utiliza una señal intermedia para saber si alguna operación del grupo DIVSQRT está en cómputo
        //assign divsqrt_busy = div_busy_o | sqrt_busy_o;

        // Generación de pulso de inicio de cada operación
        //assign div_start_i  = in_valid & ~divsqrt_busy && (op_i == fpnew_pkg::DIV);
        //assign sqrt_start_i = in_valid & ~divsqrt_busy && (op_i == fpnew_pkg::SQRT);
        
        assign lane_busy[lane]   = div_busy_o | sqrt_busy_o; // El busy está en el wrapper, aquí es 0 si está corriendo la operación.
        assign lane_in_ready[lane] = ~lane_busy[lane];


        // MUX para seleccionar las señales del módulo de DIV
        always_comb begin
          case(op_i)
            fpnew_pkg::DIV: begin
              op_result         = div_result;
              op_status         = div_status;
              out_valid         = div_out_valid;
              //lane_in_ready[lane] = in_valid & ~divsqrt_busy;
              //lane_busy[lane] = divsqrt_busy;
              //lane_in_ready[lane] = div_in_ready_o;
              //lane_busy[lane]   = div_busy_o; // El busy está en el wrapper, aquí es 0 si está corriendo la operación.
            end
            fpnew_pkg::SQRT: begin 
              op_result         = sqrt_result;
              op_status         = sqrt_status;
              out_valid         = sqrt_out_valid;
              //lane_in_ready[lane] = in_valid & ~divsqrt_busy;
              //lane_busy[lane] = divsqrt_busy;
              //lane_in_ready[lane] = sqrt_in_ready_o;
              //lane_busy[lane]   = sqrt_busy_o; // El busy está en el wrapper, aquí es 0 si está corriendo la operación.
            end
            default: begin
              op_result         = '{default: 1'bx};
              op_status         = '{default: 1'bx};
              out_valid         = 1'b0;
              //lane_in_ready[lane] = 1'b0;
              //lane_busy[lane]   = 1'b0;
            end
          endcase
        end
        assign lane_is_class[lane]   = 1'b0;
        assign lane_class_mask[lane] = fpnew_pkg::NEGINF;
        
      end else if (OpGroup == fpnew_pkg::NONCOMP) begin : lane_instance
        fpnew_noncomp #(
          .FpFormat   (FpFormat),
          .NumPipeRegs(NumPipeRegs),
          .PipeConfig (PipeConfig),
          .TagType    (TagType),
          .AuxType    (logic)
        ) i_noncomp (
          .clk_i,
          .rst_ni,
          .operands_i      ( local_operands               ),
          .is_boxed_i      ( is_boxed_i[NUM_OPERANDS-1:0] ),
          .rnd_mode_i,
          .op_i,
          .op_mod_i,
          .tag_i,
          .mask_i          ( simd_mask_i[lane]     ),
          .aux_i           ( vectorial_op          ), // Remember whether operation was vectorial
          .in_valid_i      ( in_valid              ),
          .in_ready_o      ( lane_in_ready[lane]   ),
          .flush_i,
          .result_o        ( op_result             ),
          .status_o        ( op_status             ),
          .extension_bit_o ( lane_ext_bit[lane]    ),
          .class_mask_o    ( lane_class_mask[lane] ),
          .is_class_o      ( lane_is_class[lane]   ),
          .tag_o           ( lane_tags[lane]       ),
          .mask_o          ( lane_masks[lane]      ),
          .aux_o           ( lane_vectorial[lane]  ),
          .out_valid_o     ( out_valid             ),
          .out_ready_i     ( out_ready             ),
          .busy_o          ( lane_busy[lane]       ),
          .reg_ena_i
        );
      end // ADD OTHER OPTIONS HERE

      // Handshakes are only done if the lane is actually used
      assign out_ready            = out_ready_i & ((lane == 0) | result_is_vector);
      assign lane_out_valid[lane] = out_valid   & ((lane == 0) | result_is_vector);

      // Properly NaN-box or sign-extend the slice result if not in use
      assign local_result      = (lane_out_valid[lane] | ExtRegEna) ? op_result : '{default: lane_ext_bit[0]};
      assign lane_status[lane] = (lane_out_valid[lane] | ExtRegEna) ? op_status : '0;

    // Otherwise generate constant sign-extension
    end else begin
      assign lane_out_valid[lane] = 1'b0; // unused lane
      assign lane_in_ready[lane]  = 1'b0; // unused lane
      assign local_result         = '{default: lane_ext_bit[0]}; // sign-extend/nan box
      assign lane_status[lane]    = '0;
      assign lane_busy[lane]      = 1'b0;
      assign lane_is_class[lane]  = 1'b0;
    end

    // Insert lane result into slice result
    assign slice_result[(unsigned'(lane)+1)*FP_WIDTH-1:unsigned'(lane)*FP_WIDTH] = local_result;

    // Create Classification results
    if (TrueSIMDClass && SIMD_WIDTH >= 10) begin : vectorial_true_class // true vectorial class blocks are 10bits in size
      assign slice_vec_class_result[lane*SIMD_WIDTH +: 10] = lane_class_mask[lane];
      assign slice_vec_class_result[(lane+1)*SIMD_WIDTH-1 -: SIMD_WIDTH-10] = '0;
    end else if ((lane+1)*8 <= Width) begin : vectorial_class // vectorial class blocks are 8bits in size
      assign local_sign = (lane_class_mask[lane] == fpnew_pkg::NEGINF ||
                           lane_class_mask[lane] == fpnew_pkg::NEGNORM ||
                           lane_class_mask[lane] == fpnew_pkg::NEGSUBNORM ||
                           lane_class_mask[lane] == fpnew_pkg::NEGZERO);
      // Write the current block segment
      assign slice_vec_class_result[(lane+1)*8-1:lane*8] = {
        local_sign,  // BIT 7
        ~local_sign, // BIT 6
        lane_class_mask[lane] == fpnew_pkg::QNAN, // BIT 5
        lane_class_mask[lane] == fpnew_pkg::SNAN, // BIT 4
        lane_class_mask[lane] == fpnew_pkg::POSZERO
            || lane_class_mask[lane] == fpnew_pkg::NEGZERO, // BIT 3
        lane_class_mask[lane] == fpnew_pkg::POSSUBNORM
            || lane_class_mask[lane] == fpnew_pkg::NEGSUBNORM, // BIT 2
        lane_class_mask[lane] == fpnew_pkg::POSNORM
            || lane_class_mask[lane] == fpnew_pkg::NEGNORM, // BIT 1
        lane_class_mask[lane] == fpnew_pkg::POSINF
            || lane_class_mask[lane] == fpnew_pkg::NEGINF // BIT 0
      };
    end
  end

  // ------------
  // Output Side
  // ------------
  assign result_is_vector = lane_vectorial[0];
  assign result_is_class  = lane_is_class[0];

  assign slice_regular_result = $signed({extension_bit_o, slice_result});

  localparam int unsigned CLASS_VEC_BITS = (NUM_LANES*8 > Width) ? 8 * (Width / 8) : NUM_LANES*8;

  // Pad out unused vec_class bits if each classify result is on 8 bits
  if (!(TrueSIMDClass && SIMD_WIDTH >= 10)) begin
    if (CLASS_VEC_BITS < Width) begin : pad_vectorial_class
      assign slice_vec_class_result[Width-1:CLASS_VEC_BITS] = '0;
    end
  end

  // localparam logic [Width-1:0] CLASS_VEC_MASK = 2**CLASS_VEC_BITS - 1;

  assign slice_class_result = result_is_vector ? slice_vec_class_result : lane_class_mask[0];

  // Select the proper result
  assign result_o = result_is_class ? slice_class_result : slice_regular_result;

  assign extension_bit_o                              = lane_ext_bit[0]; // upper lanes unused
  assign tag_o                                        = lane_tags[0];    // upper lanes unused
  assign busy_o                                       = (| lane_busy);
  assign out_valid_o                                  = lane_out_valid[0]; // upper lanes unused


  // Collapse the lane status
  always_comb begin : output_processing
    // Collapse the status
    automatic fpnew_pkg::status_t temp_status;
    temp_status = '0;
    for (int i = 0; i < int'(NUM_LANES); i++)
      temp_status |= lane_status[i] & {5{lane_masks[i]}};
    status_o = temp_status;
  end
endmodule
